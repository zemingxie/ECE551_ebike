package test;
  
endpackage
