module eBike_tb();
 
  // include or import tasks?

  localparam FAST_SIM = 1;		// accelerate simulation by default

  ///////////////////////////
  // Stimulus of type reg //
  /////////////////////////
  reg clk,RST_n;
  reg [11:0] BATT;				// analog values
  reg [11:0] BRAKE,TORQUE;		// analog values
  reg tgglMd;					// push button for assist mode
  reg [15:0] YAW_RT;			// models angular rate of incline (+ => uphill)


  //////////////////////////////////////////////////
  // Declare any internal signal to interconnect //
  ////////////////////////////////////////////////
  wire A2D_SS_n,A2D_MOSI,A2D_SCLK,A2D_MISO;
  wire highGrn,lowGrn,highYlw,lowYlw,highBlu,lowBlu;
  wire hallGrn,hallBlu,hallYlw;
  wire inertSS_n,inertSCLK,inertMISO,inertMOSI,inertINT;
  logic cadence;
  wire [1:0] LED;			// hook to setting from PB_intf
  
  wire signed [11:0] coilGY,coilYB,coilBG;
  logic [11:0] curr;		// comes from hub_wheel_model
  wire [11:0] BATT_TX, TORQUE_TX, CURR_TX;
  logic vld_TX;
  logic TX_RX;
  logic [7:0] rx_data;
  integer cadence_rate;
  
  //////////////////////////////////////////////////
  // Instantiate model of analog input circuitry //
  ////////////////////////////////////////////////
  AnalogModel iANLG(.clk(clk),.rst_n(RST_n),.SS_n(A2D_SS_n),.SCLK(A2D_SCLK),
                    .MISO(A2D_MISO),.MOSI(A2D_MOSI),.BATT(BATT),
		    .CURR(curr),.BRAKE(BRAKE),.TORQUE(TORQUE));

  ////////////////////////////////////////////////////////////////
  // Instantiate model inertial sensor used to measure incline //
  //////////////////////////////////////////////////////////////
  eBikePhysics iPHYS(.clk(clk),.RST_n(RST_n),.SS_n(inertSS_n),.SCLK(inertSCLK),
	             .MISO(inertMISO),.MOSI(inertMOSI),.INT(inertINT),
		     .yaw_rt(YAW_RT),.highGrn(highGrn),.lowGrn(lowGrn),
		     .highYlw(highYlw),.lowYlw(lowYlw),.highBlu(highBlu),
		     .lowBlu(lowBlu),.hallGrn(hallGrn),.hallYlw(hallYlw),
		     .hallBlu(hallBlu),.avg_curr(curr));

  //////////////////////
  // Instantiate DUT //
  ////////////////////
  eBike #(FAST_SIM) iDUT(.clk(clk),.RST_n(RST_n),.A2D_SS_n(A2D_SS_n),.A2D_MOSI(A2D_MOSI),
                         .A2D_SCLK(A2D_SCLK),.A2D_MISO(A2D_MISO),.hallGrn(hallGrn),
			 .hallYlw(hallYlw),.hallBlu(hallBlu),.highGrn(highGrn),
			 .lowGrn(lowGrn),.highYlw(highYlw),.lowYlw(lowYlw),
			 .highBlu(highBlu),.lowBlu(lowBlu),.inertSS_n(inertSS_n),
			 .inertSCLK(inertSCLK),.inertMOSI(inertMOSI),
			 .inertMISO(inertMISO),.inertINT(inertINT),
			 .cadence(cadence),.tgglMd(tgglMd),.TX(TX_RX),
			 .LED(LED));
			 
			 
  ////////////////////////////////////////////////////////////
  // Instantiate UART_rcv or some other telemetry monitor? //
  //////////////////////////////////////////////////////////
  UART_rcv ircv(.clk(clk), .rst_n(RST_n), .RX(TX_RX), .rdy(vld_TX), .rx_data(rx_data), .clr_rdy(vld_TX));
  integer prev_omega;
  integer prev_curr;
  integer prev_duty;
  integer prev_drvmag;
  initial begin
    clk = 0;
    RST_n = 0;
    TORQUE = 12'h700;
    cadence = 1'b0;
    YAW_RT = 16'h0000;
    BATT = 12'hb80;
    BRAKE = 12'hfff;
    tgglMd = 1'b0;
	cadence_rate = 2200;
    @(posedge clk);
    @(negedge clk) RST_n = 1;
	@(posedge clk);	
	repeat(500000) @(posedge clk);
	if(iDUT.error != iDUT.isensor.target_curr - iDUT.isensor.avg_curr) begin
		$display("Error is incorrect");
		$stop();
	end
	prev_omega = iPHYS.omega;
	prev_curr = iDUT.isensor.target_curr;
	repeat(500000) @(posedge clk);
	if(iDUT.error != iDUT.isensor.target_curr - iDUT.isensor.avg_curr) begin
		$display("Error is incorrect");
		$stop();
	end
	if(prev_omega >= iPHYS.omega) begin
		$display("Omega is falling when it should be rising");
	end
	if(prev_curr >= iDUT.isensor.target_curr) begin
		$display("Current is falling when it should be rising");
		$stop();
	end
	if(!(iDUT.iInert.incline == 13'h0000 || iDUT.iInert.incline == 13'h1fff)) begin
		$display("Incline is changing unexpectedly");
		$stop();
	end
	prev_duty = iDUT.ibrushless.duty;
	prev_drvmag = iDUT.iPID.drv_mag;
    	repeat(1100000) @(posedge clk);
	cadence_rate = 8192;
	TORQUE = 12'h500;
	repeat(500000) @(posedge clk);
	if(iDUT.error != iDUT.isensor.target_curr - iDUT.isensor.avg_curr) begin
		$display("Error is incorrect");
		$stop();
	end
	prev_omega = iPHYS.omega;
	prev_curr = iDUT.isensor.target_curr;
	repeat(500000) @(posedge clk);	
	if(iDUT.error != iDUT.isensor.target_curr - iDUT.isensor.avg_curr) begin
		$display("Error is incorrect");
		$stop();
	end
	if(prev_omega <= iPHYS.omega) begin
		$display("Omega is rising when it should be falling");
		$stop();
	end
	if(prev_curr <= iDUT.isensor.target_curr) begin
		$display("Current is rising when it should be falling");
		$stop();
	end
	if(!(iDUT.iInert.incline == 13'h0000 || iDUT.iInert.incline == 13'h1fff)) begin
		$display("Incline is changing unexpectedly");
		$stop();
	end
	if(iDUT.ibrushless.duty > prev_duty) begin
		$display("duty cycle higher than expected");
		$stop();
	end
	if(iDUT.iPID.drv_mag > prev_drvmag) begin
		$display("motor drive higher than expected");
		$stop();
	end
	repeat(1100000) @(posedge clk);

    $stop();
	
  end
  
  ///////////////////
  // Generate clk //
  /////////////////
  always
    #10 clk = ~clk;

  ///////////////////////////////////////////
  // Block for cadence signal generation? //
  /////////////////////////////////////////
  always begin
    repeat(cadence_rate) @(posedge clk); 
	cadence = ~cadence;		
  end
	
endmodule
