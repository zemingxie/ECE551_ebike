module cadence_LU(cadence_per,cadence);

  ///////////////////////////////////////////////////
  // Non-linear transform of cadence period to a  //
  // 5-bit vector (cadence) representing cadence //
  // Implemented in CadenceTransform.xlsx       //
  ///////////////////////////////////////////////
  input [7:0] cadence_per;
  output reg [4:0] cadence;
  
  always_comb
    case (cadence_per)
		8'h8 : cadence = 5'h1F;
		8'h9 : cadence = 5'h1F;
		8'hA : cadence = 5'h1F;
		8'hB : cadence = 5'h1F;
		8'hC : cadence = 5'h1E;
		8'hD : cadence = 5'h1D;
		8'hE : cadence = 5'h1C;
		8'hF : cadence = 5'h1B;
		8'h10 : cadence = 5'h1A;
		8'h11 : cadence = 5'h1A;
		8'h12 : cadence = 5'h19;
		8'h13 : cadence = 5'h19;
		8'h14 : cadence = 5'h18;
		8'h15 : cadence = 5'h18;
		8'h16 : cadence = 5'h17;
		8'h17 : cadence = 5'h17;
		8'h18 : cadence = 5'h17;
		8'h19 : cadence = 5'h16;
		8'h1A : cadence = 5'h16;
		8'h1B : cadence = 5'h16;
		8'h1C : cadence = 5'h16;
		8'h1D : cadence = 5'h15;
		8'h1E : cadence = 5'h15;
		8'h1F : cadence = 5'h15;
		8'h20 : cadence = 5'h15;
		8'h21 : cadence = 5'h15;
		8'h22 : cadence = 5'h14;
		8'h23 : cadence = 5'h14;
		8'h24 : cadence = 5'h14;
		8'h25 : cadence = 5'h14;
		8'h26 : cadence = 5'h14;
		8'h27 : cadence = 5'h14;
		8'h28 : cadence = 5'h13;
		8'h29 : cadence = 5'h13;
		8'h2A : cadence = 5'h13;
		8'h2B : cadence = 5'h13;
		8'h2C : cadence = 5'h13;
		8'h2D : cadence = 5'h13;
		8'h2E : cadence = 5'h13;
		8'h2F : cadence = 5'h13;
		8'h30 : cadence = 5'h13;
		8'h31 : cadence = 5'h12;
		8'h32 : cadence = 5'h12;
		8'h33 : cadence = 5'h12;
		8'h34 : cadence = 5'h12;
		8'h35 : cadence = 5'h12;
		8'h36 : cadence = 5'h12;
		8'h37 : cadence = 5'h12;
		8'h38 : cadence = 5'h12;
		8'h39 : cadence = 5'h12;
		8'h3A : cadence = 5'h12;
		8'h3B : cadence = 5'h12;
		8'h3C : cadence = 5'h12;
		8'h3D : cadence = 5'h12;
		8'h3E : cadence = 5'h12;
		8'h3F : cadence = 5'h11;
		8'h40 : cadence = 5'h11;
		8'h41 : cadence = 5'h11;
		8'h42 : cadence = 5'h11;
		8'h43 : cadence = 5'h11;
		8'h44 : cadence = 5'h11;
		8'h45 : cadence = 5'h11;
		8'h46 : cadence = 5'h11;
		8'h47 : cadence = 5'h11;
		8'h48 : cadence = 5'h11;
		8'h49 : cadence = 5'h11;
		8'h4A : cadence = 5'h11;
		8'h4B : cadence = 5'h11;
		8'h4C : cadence = 5'h11;
		8'h4D : cadence = 5'h11;
		8'h4E : cadence = 5'h11;
		8'h4F : cadence = 5'h11;
		8'h50 : cadence = 5'h11;
		8'h51 : cadence = 5'h11;
		8'h52 : cadence = 5'h11;
		8'h53 : cadence = 5'h11;
		8'h54 : cadence = 5'h11;
		8'h55 : cadence = 5'h11;
		8'h56 : cadence = 5'h11;
		8'h57 : cadence = 5'h10;
		8'h58 : cadence = 5'h10;
		8'h59 : cadence = 5'h10;
		8'h5A : cadence = 5'h10;
		8'h5B : cadence = 5'h10;
		8'h5C : cadence = 5'h10;
		8'h5D : cadence = 5'h10;
		8'h5E : cadence = 5'h10;
		8'h5F : cadence = 5'h10;
		8'h60 : cadence = 5'h10;
		8'h61 : cadence = 5'h10;
		8'h62 : cadence = 5'h10;
		8'h63 : cadence = 5'h10;
		8'h64 : cadence = 5'h10;
		8'h65 : cadence = 5'h10;
		8'h66 : cadence = 5'h10;
		8'h67 : cadence = 5'h10;
		8'h68 : cadence = 5'h10;
		8'h69 : cadence = 5'h10;
		8'h6A : cadence = 5'h10;
		8'h6B : cadence = 5'h10;
		8'h6C : cadence = 5'h10;
		8'h6D : cadence = 5'h10;
		8'h6E : cadence = 5'h10;
		8'h6F : cadence = 5'h10;
		8'h70 : cadence = 5'h10;
		8'h71 : cadence = 5'h10;
		8'h72 : cadence = 5'h10;
		8'h73 : cadence = 5'h10;
		8'h74 : cadence = 5'h10;
		8'h75 : cadence = 5'h10;
		8'h76 : cadence = 5'h10;
		8'h77 : cadence = 5'h10;
		8'h78 : cadence = 5'h10;
		8'h79 : cadence = 5'h10;
		8'h7A : cadence = 5'h10;
		8'h7B : cadence = 5'h10;
		8'h7C : cadence = 5'h10;
		8'h7D : cadence = 5'h10;
		8'h7E : cadence = 5'h10;
		8'h7F : cadence = 5'h10;
		8'h80 : cadence = 5'h10;
		8'h81 : cadence = 5'h10;
		8'h82 : cadence = 5'h10;
		8'h83 : cadence = 5'h10;
		8'h84 : cadence = 5'h10;
		8'h85 : cadence = 5'h10;
		8'h86 : cadence = 5'h10;
		8'h87 : cadence = 5'h10;
		8'h88 : cadence = 5'h10;
		8'h89 : cadence = 5'h10;
		8'h8A : cadence = 5'h10;
		8'h8B : cadence = 5'hF;
		8'h8C : cadence = 5'hF;
		8'h8D : cadence = 5'hF;
		8'h8E : cadence = 5'hF;
		8'h8F : cadence = 5'hF;
		8'h90 : cadence = 5'hF;
		8'h91 : cadence = 5'hF;
		8'h92 : cadence = 5'hF;
		8'h93 : cadence = 5'hF;
		8'h94 : cadence = 5'hF;
		8'h95 : cadence = 5'hF;
		8'h96 : cadence = 5'hF;
		8'h97 : cadence = 5'hF;
		8'h98 : cadence = 5'hF;
		8'h99 : cadence = 5'hF;
		8'h9A : cadence = 5'hF;
		8'h9B : cadence = 5'hF;
		8'h9C : cadence = 5'hF;
		8'h9D : cadence = 5'hF;
		8'h9E : cadence = 5'hF;
		8'h9F : cadence = 5'hF;
		8'hA0 : cadence = 5'hF;
		8'hA1 : cadence = 5'hF;
		8'hA2 : cadence = 5'hF;
		8'hA3 : cadence = 5'hF;
		8'hA4 : cadence = 5'hF;
		8'hA5 : cadence = 5'hF;
		8'hA6 : cadence = 5'hF;
		8'hA7 : cadence = 5'hF;
		8'hA8 : cadence = 5'hF;
		8'hA9 : cadence = 5'hF;
		8'hAA : cadence = 5'hF;
		8'hAB : cadence = 5'hF;
		8'hAC : cadence = 5'hF;
		8'hAD : cadence = 5'hF;
		8'hAE : cadence = 5'hF;
		8'hAF : cadence = 5'hF;
		8'hB0 : cadence = 5'hF;
		8'hB1 : cadence = 5'hF;
		8'hB2 : cadence = 5'hF;
		8'hB3 : cadence = 5'hF;
		8'hB4 : cadence = 5'hF;
		8'hB5 : cadence = 5'hF;
		8'hB6 : cadence = 5'hF;
		8'hB7 : cadence = 5'hF;
		8'hB8 : cadence = 5'hF;
		8'hB9 : cadence = 5'hF;
		8'hBA : cadence = 5'hF;
		8'hBB : cadence = 5'hF;
		8'hBC : cadence = 5'hF;
		8'hBD : cadence = 5'hF;
		8'hBE : cadence = 5'hF;
		8'hBF : cadence = 5'hF;
		8'hC0 : cadence = 5'hF;
		8'hC1 : cadence = 5'hF;
		8'hC2 : cadence = 5'hF;
		8'hC3 : cadence = 5'hF;
		8'hC4 : cadence = 5'hF;
		8'hC5 : cadence = 5'hF;
		8'hC6 : cadence = 5'hF;
		8'hC7 : cadence = 5'hF;
		8'hC8 : cadence = 5'hF;
		8'hC9 : cadence = 5'hF;
		8'hCA : cadence = 5'hF;
		8'hCB : cadence = 5'hF;
		8'hCC : cadence = 5'hF;
		8'hCD : cadence = 5'hF;
		8'hCE : cadence = 5'hF;
		8'hCF : cadence = 5'hF;
		8'hD0 : cadence = 5'hF;
		8'hD1 : cadence = 5'hF;
		8'hD2 : cadence = 5'hF;
		8'hD3 : cadence = 5'hF;
		8'hD4 : cadence = 5'hF;
		8'hD5 : cadence = 5'hF;
		8'hD6 : cadence = 5'hF;
		8'hD7 : cadence = 5'hF;
		8'hD8 : cadence = 5'hF;
		8'hD9 : cadence = 5'hF;
		8'hDA : cadence = 5'hF;
		8'hDB : cadence = 5'hF;
		8'hDC : cadence = 5'hF;
		8'hDD : cadence = 5'hF;
		8'hDE : cadence = 5'hF;
		8'hDF : cadence = 5'hF;
		8'hE0 : cadence = 5'hF;
		8'hE1 : cadence = 5'hF;
		8'hE2 : cadence = 5'hF;
		8'hE3 : cadence = 5'hF;
		8'hE4 : cadence = 5'hF;
		default : cadence = 5'hF;
	endcase

endmodule